----------------------------------------------------------------------------------
-- Archivo autogenerado con 'converter.cpp'
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

use work.tipos.all;

entity vga_RecButton is
	generic(N: integer := 62; M: integer := 13);
	port(
		hcnt: in std_logic_vector(8 downto 0);
		vcnt: in std_logic_vector(9 downto 0);
		hcnt_aux: in std_logic_vector(8 downto 0);
		vcnt_aux: in std_logic_vector(9 downto 0);
		pintar: out std_logic;
		currentobject: out vga_object --el tipo vga_object esta definido en tipos.vhd
	);
end vga_recButton;

architecture arch of vga_RecButton is

type vga_RecButton_img_type is array (M*2 - 1 downto 0) of std_logic_vector(N - 1 downto 0);
signal vga_RecButton_img : vga_RecButton_img_type := (
"00011111110000000111111100001111111111000111110000000000000000", "00011111110000000111111100001111111111000111110000000000000000", 
"00111111111000000111111110001111111111001111111100000000000000", "00111111111000000111111110001111111111001111111100000000000000", 
"01111111111100000110000011101100000000011100001110000000000000", "01111111111100000110000011101100000000011100001110000000000000", 
"11111111111110000110000011101100000000011000001110000000000000", "11111111111110000110000011101100000000011000001110000000000000", 
"11111111111110000110000011101100000000011000000000000000000000", "11111111111110000110000011101100000000011000000000000000000000", 
"11111111111110000110000011101111111100011000000000000000000000", "11111111111110000110000011101111111100011000000000000000000000", 
"11111111111110000111111111101111111100011000000000000000000000", "11111111111110000111111111101111111100011000000000000000000000", 
"11111111111110000111111111001100000000011000000000000000000000", "11111111111110000111111111001100000000011000000000000000000000", 
"11111111111110000111111110001100000000011000000000000000000000", "11111111111110000111111110001100000000011000000000000000000000", 
"11111111111110000110000111001100000000011000001110000000000000", "11111111111110000110000111001100000000011000001110000000000000", 
"01111111111100000110000011101100000000011100001110000000000000", "01111111111100000110000011101100000000011100001110000000000000", 
"00111111111000000110000011101111111111011111111110000000000000", "00111111111000000110000011101111111111011111111110000000000000", 
"00011111110000000110000011101111111111001111111000000000000000", "00011111110000000110000011101111111111001111111000000000000000");

begin

currentobject <= teclaPulsada; --Modificar el objeto para el color que se necesite

pintar_vga_RecButton: process(hcnt, vcnt)
begin
	if hcnt - hcnt_aux > N-1 or vcnt - vcnt_aux > M*2 - 1 then
		pintar <= '0';
	else pintar <= vga_RecButton_img(conv_integer(M*2 - 1 - vcnt + vcnt_aux))(conv_integer(N - 1 - hcnt + hcnt_aux));
	end if;

end process;

end arch;

