----------------------------------------------------------------------------------
-- Archivo autogenerado con 'converter.cpp'
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

use work.tipos.all;

entity vga_playButton is
	generic(N: integer := 62; M: integer := 13);
	port(
		hcnt: in std_logic_vector(8 downto 0);
		vcnt: in std_logic_vector(9 downto 0);
		hcnt_aux: in std_logic_vector(8 downto 0);
		vcnt_aux: in std_logic_vector(9 downto 0);
		pintar: out std_logic;
		currentobject: out vga_object --el tipo vga_object esta definido en tipos.vhd
	);
end vga_playButton;

architecture arch of vga_playButton is

type vga_playButton_img_type is array (M*2 - 1 downto 0) of std_logic_vector(N - 1 downto 0);
signal vga_playButton_img : vga_playButton_img_type := (
"11110000000000001111111100111000000000011111100011000001110000", "11110000000000001111111100111000000000011111100011000001110000", 
"11111100000000001111111100111000000000011111100011000001110000", "11111100000000001111111100111000000000011111100011000001110000", 
"11111111000000001100000110111000000001110000111011000001110000", "11111111000000001100000110111000000001110000111011000001110000", 
"11111111110000001100000110111000000001110000111011110111110000", "11111111110000001100000110111000000001110000111011110111110000", 
"11111111111100001100000110111000000001110000111000110111000000", "11111111111100001100000110111000000001110000111000110111000000", 
"11111111111110001100000110111000000001110000111000111111000000", "11111111111110001100000110111000000001110000111000111111000000", 
"11111111111111001111111110111000000001111111111000111111000000", "11111111111111001111111110111000000001111111111000111111000000", 
"11111111111110001111111100111000000001111111111000011100000000", "11111111111110001111111100111000000001111111111000011100000000", 
"11111111111100001111111000111000000001111111111000011100000000", "11111111111100001111111000111000000001111111111000011100000000", 
"11111111110000001100000000111000000001110000111000011100000000", "11111111110000001100000000111000000001110000111000011100000000", 
"11111111000000001100000000111000000001110000111000011100000000", "11111111000000001100000000111000000001110000111000011100000000", 
"11111100000000001100000000111111111101110000111000011100000000", "11111100000000001100000000111111111101110000111000011100000000", 
"11110000000000001100000000111111111101110000111000011100000000", "11110000000000001100000000111111111101110000111000011100000000");

begin

currentobject <= colorVerde; --Modificar el objeto para el color que se necesite

pintar_vga_playButton: process(hcnt, vcnt)
begin
	if hcnt - hcnt_aux > N or vcnt - vcnt_aux > M*2 then
		pintar <= '0';
	else pintar <= vga_playButton_img(conv_integer(M*2 - 1 - vcnt + vcnt_aux))(conv_integer(N - 1 - hcnt + hcnt_aux));
	end if;

end process;

end arch;