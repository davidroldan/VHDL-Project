----------------------------------------------------------------------------------
-- Archivo autogenerado con 'converter.cpp'
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

use work.tipos.all;

entity vga_stopButton is
	generic(N: integer := 62; M: integer := 13);
	port(
		hcnt: in std_logic_vector(8 downto 0);
		vcnt: in std_logic_vector(9 downto 0);
		hcnt_aux: in std_logic_vector(8 downto 0);
		vcnt_aux: in std_logic_vector(9 downto 0);
		pintar: out std_logic;
		currentobject: out vga_object --el tipo vga_object esta definido en tipos.vhd
	);
end vga_stopButton;

architecture arch of vga_stopButton is

type vga_stopButton_img_type is array (M*2 - 1 downto 0) of std_logic_vector(N - 1 downto 0);
signal vga_stopButton_img : vga_stopButton_img_type := (
"11111111111110000111111100111111111100011111100001111111100000", "11111111111110000111111100111111111100011111100001111111100000", 
"11111111111110001111111100111111111100111111110001111111110000", "11111111111110001111111100111111111100111111110001111111110000", 
"11111111111110001110000000111111111100111001110001110001111000", "11111111111110001110000000111111111100111001110001110001111000", 
"11111111111110001100000000000111100000111001110001110000111000", "11111111111110001100000000000111100000111001110001110000111000", 
"11111111111110001110000000000111100001111001111001110001111000", "11111111111110001110000000000111100001111001111001110001111000", 
"11111111111110001111111100000111100001111001111001111111111000", "11111111111110001111111100000111100001111001111001111111111000", 
"11111111111110000111111110000111100001111001111001111111110000", "11111111111110000111111110000111100001111001111001111111110000", 
"11111111111110000000001110000111100001111001111001111111100000", "11111111111110000000001110000111100001111001111001111111100000", 
"11111111111110000000001110000111100001111001111001110000000000", "11111111111110000000001110000111100001111001111001110000000000", 
"11111111111110000000001110000111100001111001111001110000000000", "11111111111110000000001110000111100001111001111001110000000000", 
"11111111111110001111111110000111100000111001110001110000000000", "11111111111110001111111110000111100000111001110001110000000000", 
"11111111111110001111111100000111100000111111110001110000000000", "11111111111110001111111100000111100000111111110001110000000000", 
"11111111111110001111111000000111100000011111100001110000000000", "11111111111110001111111000000111100000011111100001110000000000");

begin

currentobject <= colorAmarillo; --Modificar el objeto para el color que se necesite

pintar_vga_stopButton: process(hcnt, vcnt)
begin
	if hcnt - hcnt_aux > N - 1 or vcnt - vcnt_aux > M*2 - 1 then
		pintar <= '0';
	else pintar <= vga_stopButton_img(conv_integer(M*2 - 1 - vcnt + vcnt_aux))(conv_integer(N - 1 - hcnt + hcnt_aux));
	end if;

end process;

end arch;